`timescale 1ns / 1ps
`include "SKELETON.v"

module tb_SKELETON();
endmodule
