//Verilog HDL for "DIGITAL", "SKELETON", "functional"


module SKELETON ();
endmodule
