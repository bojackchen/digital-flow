`timescale 1ns / 1ps
`include "SKELETON_syn.v"

module tb_SKELETON();
endmodule
