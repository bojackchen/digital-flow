`timescale 1ns / 1ps
`include "SKELETON_encounter.v"

module tb_SKELETON();
endmodule
